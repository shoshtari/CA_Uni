Add d0, d1
Add d0, 25
Subtract d0, d1
Addi d0, 50
And d0, d1
Sll d0, 10
Lw d0, 7
Sw d0, 10
CLR d0
Mov BA, 50
CMP d0, d1
Bne 25
Jmp 2500